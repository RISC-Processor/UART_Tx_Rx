module DataMemWrapper (
	input logic  clk,
	input logic  rst
);




endmodule